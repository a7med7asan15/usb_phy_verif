//  Interface: usbf_intf
//
interface utmi_intf(input clk, reset);

    
endinterface: utmi_intf
