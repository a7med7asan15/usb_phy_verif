package env_pkg;
    import uvm_pkg::*;
    `include "uvm_macros.svh"

    import top_params_pkg::*;
    import riscv_pkg::*; 

    `include "src/d_env_config.svh"
    `include "src/d_env.svh"
    
endpackage: env_pkg
