package seq_pkg;
    import uvm_pkg::*;
    `include "uvm_macros.svh"
    
    import top_params_pkg::*;

    `include "src/riscv_sequence_items/riscv_seq_item.svh"
    `include "src/riscv_sequence_items/b_seq_item.svh"
    `include "src/riscv_sequence_items/i_seq_item.svh"
    `include "src/riscv_sequence_items/j_seq_item.svh"
    `include "src/riscv_sequence_items/s_seq_item.svh"
    `include "src/riscv_sequence_items/u_seq_item.svh"
    `include "src/riscv_sequence_items/r_seq_item.svh"
    `include "src/riscv_sequences/base_sequence.svh"
    `include "src/riscv_sequences/random_sequence.svh"
    `include "src/riscv_sequencer.svh"

endpackage: seq_pkg
