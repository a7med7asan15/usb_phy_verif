//  Interface: usbf_intf
//
interface sram_intf
    /*  package imports  */
    #(
        <parameter_list>
    )(
        <port_list>
    );

    
endinterface: sram_intf
