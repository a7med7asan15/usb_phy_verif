//  Interface: usbf_intf
//
interface usbf_intf
    /*  package imports  */
    #(
        <parameter_list>
    )(
        <port_list>
    );

    
endinterface: usbf_intf
