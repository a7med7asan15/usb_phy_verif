package analysis_pkg;
    import uvm_pkg::*;
    `include "uvm_macros.svh"

    import top_params_pkg::*;
    import seq_pkg::*;

    `include "src/riscv_scoreboard.svh"
    `include "src/riscv_subscriber.svh"
    
endpackage: analysis_pkg
