package top_params_pkg;


endpackage: top_params_pkg